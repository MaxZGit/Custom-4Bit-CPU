`timescale 10ns/1ps


`include "src/half_adder.v"
`include "src/full_adder.v"
`include "src/carry_ripple_adder.v"
`include "src/alu.v"
`include "src/my_register.v"
`include "src/reg_memory.v"
`include "src/control_unit.v"
`include "src/cpu.v"
`include "src/uart_rx.v"
`include "src/programmer.v"


module cpu_tb;
    
    // Instruction constants
    localparam NOP_INSTR = 4'b0000;
    localparam XOR_INSTR = 4'b0001;
    localparam AND_INSTR = 4'b0010;
    localparam OR_INSTR = 4'b0011;
    localparam ADD_INSTR = 4'b0100;
    localparam INC_INSTR = 4'b0101;
    localparam DEC_INSTR = 4'b0110;
    localparam SUB_INSTR = 4'b0111;
    localparam JMP_INSTR = 4'b1000;
    localparam JZ_INSTR = 4'b1001;
    localparam JC_INSTR = 4'b1010;
    localparam LD_INSTR = 4'b1011;
    localparam ST_INSTR = 4'b1100;
    localparam IN_INSTR = 4'b1101;
    localparam OUT_INSTR = 4'b1110;
    localparam LDI_INSTR = 4'b1111;

    // ---------------------------------
    // Test programs
    // ---------------------------------

    // _._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._
    // expected behaviour: 
    // out_pins => 0001 -> 0010 -> 0100 -> 1000 -> 0001 ...
    // _._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._
    localparam TEST_CIRC_LEFT_SHIFT = 0;
    reg [63:0] circ_left_shift;  // holds 8 bytes (8 × 8 bits)
    initial begin
        circ_left_shift = {
            IN_INSTR,          // A <- IN
            OUT_INSTR,         // OUT <- A
            ST_INSTR,  4'b1111,// MEM[15] <- A
            ADD_INSTR, 4'b1111,// A <- A + MEM[15]
            JC_INSTR,  4'b1010,// if carry: jump
            JMP_INSTR, 4'b0001,// jump to OUT
            INC_INSTR,         // A <- A + 1
            JMP_INSTR, 4'b0001, // jump to OUT
            NOP_INSTR,
            NOP_INSTR,
            4'b0001
        };
    end

    // _._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._
    // expected behaviour:
    // out_pins => 0000 -> 0001 -> 0010 -> 0011 -> 0100 -> ...
    // _._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._

    localparam TEST_INC_COUNTER = 1;
    reg [63:0] inc_counter;

    initial begin
        inc_counter = {
            LDI_INSTR, 4'b0000,// A <- 0
            OUT_INSTR,         // OUT <- A
            INC_INSTR,         // A <- A + 1
            JMP_INSTR, 4'b0001,// loop back to OUT
            NOP_INSTR,
            NOP_INSTR,
            NOP_INSTR,
            NOP_INSTR,
            NOP_INSTR,
            NOP_INSTR,
            NOP_INSTR,
            NOP_INSTR,
            NOP_INSTR,
            NOP_INSTR
        };
    end

    // _._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._
    // expected behaviour:
    // out_pins: 0000 -> 1111 -> 0000 -> 1111 ...
    // _._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._

    localparam TEST_BLINK = 2;
    reg [63:0] blink;

    initial begin
        blink = {
            LDI_INSTR, 4'b0000, 
            OUT_INSTR,          
            LDI_INSTR, 4'b1111,
            OUT_INSTR,
            JMP_INSTR,  4'b0000

        };
    end

    // _._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._
    // expected behaviour:
    // out_pins => 1010 (value stored and reloaded from memory)
    // tests ST and LD instructions
    // _._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._

    localparam TEST_MEM_RW = 3;
    reg [63:0] mem_rw_test;

    initial begin
        mem_rw_test = {
            LDI_INSTR, 4'b1010,// A <- 10
            ST_INSTR,  4'b0011,// MEM[3] <- A
            LDI_INSTR, 4'b0000,// A <- 0
            LD_INSTR,  4'b0011,// A <- MEM[3]
            OUT_INSTR,         // OUT <- A
            JMP_INSTR, 4'b0100,// loop at OUT
            NOP_INSTR,
            NOP_INSTR,
            NOP_INSTR,
            NOP_INSTR,
            NOP_INSTR
        };
    end

    
    // _._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._
    // LED effect: input mirror
    // expected behaviour: LEDs follow input
    // _._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._._

    localparam TEST_INPUT_ECHO = 4;
    reg [63:0] input_echo;

    initial begin
        input_echo = {
            IN_INSTR,           // A <- IN
            OUT_INSTR,          // OUT <- A
            JMP_INSTR, 4'b0000, // loop
            NOP_INSTR,
            NOP_INSTR,
            NOP_INSTR,
            NOP_INSTR,
            NOP_INSTR
        };
    end

    localparam OPERATION_CODE_WIDTH = 3;
    localparam CRA_BIT_NUMB = 4;
    localparam REGISTER_WIDTH = 4;
    localparam MEMORY_ADDRESS_WIDTH = 4;
    localparam MEMORY_REGISTERS = 16;

    localparam UART_DATA_LENGTH = 8;
    localparam RX_COUNTER_BITWIDTH = 3;
    localparam BAUD_COUNTS_PER_BIT = 521; // for 10MHz clk
    localparam BAUD_RATE_COUNTER_BITWIDTH = 10; //2^10 0 1024
    
    localparam clk_pulse = 10;
    localparam wait_one_bit = 10*521;
    integer i;
    integer j;

    reg reset_tb = 1'b1;
    reg clk_tb = 1'b1;
    reg [REGISTER_WIDTH - 1:0] in_pins_tb = 4'b0010;
    wire [REGISTER_WIDTH - 1:0] out_pins_tb;

    reg p_program_tb = 0;
    reg rx_tb = 1;

    reg [63:0] data_array;  // holds 8 bytes (8 × 8 bits)
    reg [7:0] current_byte;

    wire next_data_strb_tb;
    wire data_valid_strb_tb;
    wire program_o_tb;
    wire fetch_instr_tb;
    wire decode_tb;
    wire fetcho_op_tb;
    wire fetch_mdr_tb;
    wire execute_tb;

    // ------------------------------------------
    // SELECT TEST PROGRAM
    // ------------------------------------------

    localparam SELECTED_TEST = TEST_INPUT_ECHO;
    
    always @(*) begin
        case (SELECTED_TEST)
            TEST_CIRC_LEFT_SHIFT: data_array = circ_left_shift;
            TEST_INC_COUNTER:     data_array = inc_counter;
            TEST_BLINK:             data_array = blink;
            TEST_MEM_RW:          data_array = mem_rw_test;
            TEST_INPUT_ECHO:          data_array = input_echo;
            default:             data_array = 64'b0;
        endcase
    end

    cpu #(
        .CRA_BIT_NUMB(CRA_BIT_NUMB),
        .OPERATION_CODE_WIDTH(OPERATION_CODE_WIDTH),
        .REGISTER_WIDTH(REGISTER_WIDTH),
        .MEMORY_ADDRESS_WIDTH(MEMORY_ADDRESS_WIDTH),
        .MEMORY_REGISTERS(MEMORY_REGISTERS),

        .UART_DATA_LENGTH(UART_DATA_LENGTH),
        .RX_COUNTER_BITWIDTH(RX_COUNTER_BITWIDTH),
        .BAUD_COUNTS_PER_BIT(BAUD_COUNTS_PER_BIT),
        .BAUD_RATE_COUNTER_BITWIDTH(BAUD_RATE_COUNTER_BITWIDTH)
    ) dut (
        .clk_i(clk_tb),
        .reset_i(reset_tb),

        .in_pins_i(in_pins_tb),
        .next_data_strb_o(next_data_strb_tb),

        .out_pins_o(out_pins_tb),
        .data_valid_strb_o(data_valid_strb_tb),

        // Status Flags
        .program_o(program_o_tb),
        .fetch_instr_o(fetch_instr_tb),
        .decode_o(decode_tb),
        .fetcho_op_o(fetcho_op_tb),
        .fetch_mdr_o(fetch_mdr_tb),
        .execute_o(execute_tb),

        .p_program_i(p_program_tb),
        .rx_i(rx_tb)
    );

    initial begin
        forever #5 clk_tb = ~clk_tb;    // Toggle clock every 5 time units
    end

    initial begin

        $dumpfile("sim/cpu_tb.vcd");
		$dumpvars;

        for (i = 0; i < MEMORY_REGISTERS; i = i + 1) begin
            $dumpvars(1, dut.memory.reg_vals[i]); // dump each element separately
        end

        reset_tb = 1'b1; // reset
        #(10*clk_pulse);
        reset_tb = 0; //release reset
        #(10*clk_pulse);

        #(1000*clk_pulse);

        p_program_tb = 1;
        for (i = 7; i >= 0; i = i - 1) begin
            current_byte = data_array[i*8+: 8];
            //start bit
            rx_tb = 0;
            #wait_one_bit;

            for (j = 0; j < 8; j = j+1) begin
                rx_tb = current_byte[j];
                #wait_one_bit;
            end

            // stop bot
            rx_tb = 1;
            #wait_one_bit;
        end

        rx_tb = 1;
        #(5*clk_pulse);
        p_program_tb = 0;

        #(1000*clk_pulse);

        $finish;
    end
endmodule